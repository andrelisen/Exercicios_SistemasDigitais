library verilog;
use verilog.vl_types.all;
entity PO_Sub_vlg_vec_tst is
end PO_Sub_vlg_vec_tst;
